-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Sun Oct 29 15:42:16 2023

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY PRUEBA IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        S_D : IN STD_LOGIC := '0';
        S_I : IN STD_LOGIC := '0';
        S : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
    );
END PRUEBA;

ARCHITECTURE BEHAVIOR OF PRUEBA IS
    TYPE type_fstate IS (state1,state2,state3);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,S_D,S_I)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= state1;
            S <= "000";
        ELSE
            S <= "000";
            CASE fstate IS
                WHEN state1 =>
                    IF (((S_D = '0') AND (S_I = '1'))) THEN
                        reg_fstate <= state1;
                    ELSE
                        reg_fstate <= state2;
                    END IF;

                    S <= "111";
                WHEN state2 =>
                    IF (((S_D = '0') AND (S_I = '1'))) THEN
                        reg_fstate <= state3;
                    ELSE
                        reg_fstate <= state2;
                    END IF;

                    S <= "101";
                WHEN state3 =>
                    IF (((S_D = '0') AND (S_I = '1'))) THEN
                        reg_fstate <= state1;
                    ELSE
                        reg_fstate <= state3;
                    END IF;

                    S <= "000";
                WHEN OTHERS => 
                    S <= "XXX";
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
