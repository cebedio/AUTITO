-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Mon Oct 23 12:14:32 2023

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY counter_16 IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        x : IN STD_LOGIC := '0';
        Z : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
    );
END counter_16;

ARCHITECTURE BEHAVIOR OF counter_16 IS
    TYPE type_fstate IS (state1,state2,state3,state4,state5,state6,state7,state8,state9,state10,state11,state12,state13,state14,state15,state16);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,x)
    BEGIN
        IF (reset='0') THEN
            reg_fstate <= state1;
            Z <= "0000";
        ELSE
            Z <= "0000";
            CASE fstate IS
                WHEN state1 =>
                    IF ((x = '1')) THEN
                        reg_fstate <= state2;
                    ELSIF ((x = '0')) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state1;
                    END IF;

                    Z <= "0000";
                WHEN state2 =>
                    IF ((x = '1')) THEN
                        reg_fstate <= state3;
                    ELSIF ((x = '0')) THEN
                        reg_fstate <= state2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state2;
                    END IF;

                    Z <= "0001";
                WHEN state3 =>
                    IF ((x = '1')) THEN
                        reg_fstate <= state4;
                    ELSIF ((x = '0')) THEN
                        reg_fstate <= state3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state3;
                    END IF;

                    Z <= "0010";
                WHEN state4 =>
                    IF ((x = '1')) THEN
                        reg_fstate <= state5;
                    ELSIF ((x = '0')) THEN
                        reg_fstate <= state4;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state4;
                    END IF;

                    Z <= "0011";
                WHEN state5 =>
                    IF ((x = '1')) THEN
                        reg_fstate <= state6;
                    ELSIF ((x = '0')) THEN
                        reg_fstate <= state5;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state5;
                    END IF;

                    Z <= "0100";
                WHEN state6 =>
                    IF ((x = '1')) THEN
                        reg_fstate <= state7;
                    ELSIF ((x = '0')) THEN
                        reg_fstate <= state6;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state6;
                    END IF;

                    Z <= "0101";
                WHEN state7 =>
                    IF ((x = '1')) THEN
                        reg_fstate <= state8;
                    ELSIF ((x = '0')) THEN
                        reg_fstate <= state7;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state7;
                    END IF;

                    Z <= "0110";
                WHEN state8 =>
                    IF ((x = '1')) THEN
                        reg_fstate <= state9;
                    ELSIF ((x = '0')) THEN
                        reg_fstate <= state8;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state8;
                    END IF;

                    Z <= "0111";
                WHEN state9 =>
                    IF ((x = '1')) THEN
                        reg_fstate <= state10;
                    ELSIF ((x = '0')) THEN
                        reg_fstate <= state9;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state9;
                    END IF;

                    Z <= "1000";
                WHEN state10 =>
                    IF ((x = '1')) THEN
                        reg_fstate <= state11;
                    ELSIF ((x = '0')) THEN
                        reg_fstate <= state10;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state10;
                    END IF;

                    Z <= "1001";
                WHEN state11 =>
                    IF ((x = '1')) THEN
                        reg_fstate <= state12;
                    ELSIF ((x = '0')) THEN
                        reg_fstate <= state11;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state11;
                    END IF;

                    Z <= "1010";
                WHEN state12 =>
                    IF ((x = '1')) THEN
                        reg_fstate <= state13;
                    ELSIF ((x = '0')) THEN
                        reg_fstate <= state12;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state12;
                    END IF;

                    Z <= "1011";
                WHEN state13 =>
                    IF ((x = '1')) THEN
                        reg_fstate <= state14;
                    ELSIF ((x = '0')) THEN
                        reg_fstate <= state13;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state13;
                    END IF;

                    Z <= "1100";
                WHEN state14 =>
                    IF ((x = '1')) THEN
                        reg_fstate <= state15;
                    ELSIF ((x = '0')) THEN
                        reg_fstate <= state14;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state14;
                    END IF;

                    Z <= "1101";
                WHEN state15 =>
                    IF ((x = '1')) THEN
                        reg_fstate <= state16;
                    ELSIF ((x = '0')) THEN
                        reg_fstate <= state15;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state15;
                    END IF;

                    Z <= "1110";
                WHEN state16 =>
                    IF ((x = '1')) THEN
                        reg_fstate <= state1;
                    ELSIF ((x = '0')) THEN
                        reg_fstate <= state16;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state16;
                    END IF;

                    Z <= "1111";
                WHEN OTHERS => 
                    Z <= "XXXX";
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
