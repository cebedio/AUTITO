library verilog;
use verilog.vl_types.all;
entity autito_principal_vlg_vec_tst is
end autito_principal_vlg_vec_tst;
